`include "bpb.vh"

/**
 * ENTRIES          : number of entries in the branch predictor buffer
 * TAG_WIDTH        : index bits
 * instr_adr        : if this address has been recorded, then CPU can go as the BPB directs
 * isbranch         : in order to register the branch when first meeted
 * real_taken       : whether this branch should be taken according to the semantics of the instructions
 * real_adr         : where should this branch jumps to
 * predict_taken    : whether this branch should be taken according to the prediction of our BPB
 * predict_adr      : where should this branch jumps to if it's taken
 */
module bpb #(
    parameter ENTRIES = `BPB_E,
    parameter TAG_WIDTH = `BPB_T
) (
    input logic clk, reset, stall, flush,
    input logic [TAG_WIDTH-1:0] instr_adr,
    input logic isbranch,
    // reality
    input logic real_taken,
    input [31:0] real_adr,
    // prediction
    output reg              predict_taken,
    output reg [31:0]       predict_adr
);

/**
 * TODO: Your code here
 */

endmodule